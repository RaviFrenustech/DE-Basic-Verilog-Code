module mux4 (
    input [1:0] sel,
    input [7:0] a,b,c,d,
    input [7:0] y
);

endmodule