module xor2 ( m1, m2, o1);

input m1, m2;
output o1;

assign o1 = m1 ^ m2;

endmodule